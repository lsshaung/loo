/*--------------------------------------
// AXI PKG
// file : axi_seq_lib_pkg.sv
// author : SeanChen
// date : 2013/05/06
// notes
---------------------------------------*/

`ifndef AXI_SEQ_LIB_PKG_SV
`define AXI_SEQ_LIB_PKG_SV

`include "../tc/testcase/sequence_libs/axi_based_seq_lib.sv"
`include "../tc/testcase/sequence_libs/axi_master_seq_lib.sv"
`include "../tc/testcase/sequence_libs/axi_master_based_seq_lib.sv"
`include "../tc/testcase/sequence_libs/axi_slave_based_seq_lib.sv"

`endif  // AXI_SEQ_LIB_PKG_SV
